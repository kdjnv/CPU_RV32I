// Created with Corsair v1.0.4

`ifndef __REGS_I2C_VH
`define __REGS_I2C_VH

`define I2C_BASE_ADDR 0
`define I2C_DATA_WIDTH 32
`define I2C_ADDR_WIDTH 32

// I2C_CONTROL - I2C Control Register
`define I2C_I2C_CONTROL_ADDR 32'h0
`define I2C_I2C_CONTROL_RESET 32'h2880a50e

// I2C_CONTROL.CLKDIV - Clock divider for SCL
`define I2C_I2C_CONTROL_CLKDIV_WIDTH 10
`define I2C_I2C_CONTROL_CLKDIV_LSB 0
`define I2C_I2C_CONTROL_CLKDIV_MASK 32'h0
`define I2C_I2C_CONTROL_CLKDIV_RESET 10'h10e

// I2C_CONTROL.NUMBRX - Number of bytes to receive (0 means 1)
`define I2C_I2C_CONTROL_NUMBRX_WIDTH 3
`define I2C_I2C_CONTROL_NUMBRX_LSB 10
`define I2C_I2C_CONTROL_NUMBRX_MASK 32'h0
`define I2C_I2C_CONTROL_NUMBRX_RESET 3'h1

// I2C_CONTROL.DUTYSCL - Duty cycle for SCL (reserved for future use)
`define I2C_I2C_CONTROL_DUTYSCL_WIDTH 4
`define I2C_I2C_CONTROL_DUTYSCL_LSB 13
`define I2C_I2C_CONTROL_DUTYSCL_MASK 32'h0
`define I2C_I2C_CONTROL_DUTYSCL_RESET 4'h5

// I2C_CONTROL.RSE - Register Slave Enable
`define I2C_I2C_CONTROL_RSE_WIDTH 1
`define I2C_I2C_CONTROL_RSE_LSB 17
`define I2C_I2C_CONTROL_RSE_MASK 32'h0
`define I2C_I2C_CONTROL_RSE_RESET 1'h0

// I2C_CONTROL.LENADD - Slave address length
`define I2C_I2C_CONTROL_LENADD_WIDTH 2
`define I2C_I2C_CONTROL_LENADD_LSB 18
`define I2C_I2C_CONTROL_LENADD_MASK 32'h0
`define I2C_I2C_CONTROL_LENADD_RESET 2'h0

// I2C_CONTROL.EN - Enable I2C
`define I2C_I2C_CONTROL_EN_WIDTH 1
`define I2C_I2C_CONTROL_EN_LSB 20
`define I2C_I2C_CONTROL_EN_MASK 32'h0
`define I2C_I2C_CONTROL_EN_RESET 1'h0

// I2C_CONTROL.STRX - Start transmit/receive
`define I2C_I2C_CONTROL_STRX_WIDTH 1
`define I2C_I2C_CONTROL_STRX_LSB 21
`define I2C_I2C_CONTROL_STRX_MASK 32'h0
`define I2C_I2C_CONTROL_STRX_RESET 1'h0

// I2C_CONTROL.MODE - Transfer mode (0 transmit, 1 receive)
`define I2C_I2C_CONTROL_MODE_WIDTH 1
`define I2C_I2C_CONTROL_MODE_LSB 22
`define I2C_I2C_CONTROL_MODE_MASK 32'h0
`define I2C_I2C_CONTROL_MODE_RESET 1'h0

// I2C_CONTROL.NUMBTX - Number of bytes to transmit (0 means 1)
`define I2C_I2C_CONTROL_NUMBTX_WIDTH 3
`define I2C_I2C_CONTROL_NUMBTX_LSB 23
`define I2C_I2C_CONTROL_NUMBTX_MASK 32'h0
`define I2C_I2C_CONTROL_NUMBTX_RESET 3'h1

// I2C_CONTROL.RST - Repeat start condition
`define I2C_I2C_CONTROL_RST_WIDTH 1
`define I2C_I2C_CONTROL_RST_LSB 26
`define I2C_I2C_CONTROL_RST_MASK 32'h0
`define I2C_I2C_CONTROL_RST_RESET 1'h0

// I2C_CONTROL.SEML - Sample location on SCL pulse (max 9)
`define I2C_I2C_CONTROL_SEML_WIDTH 5
`define I2C_I2C_CONTROL_SEML_LSB 27
`define I2C_I2C_CONTROL_SEML_MASK 32'h0
`define I2C_I2C_CONTROL_SEML_RESET 5'h5


// I2C_STATUS - I2C Status Register
`define I2C_I2C_STATUS_ADDR 32'h4
`define I2C_I2C_STATUS_RESET 32'h42

// I2C_STATUS.SLAVE_FOUND - Slave address detected
`define I2C_I2C_STATUS_SLAVE_FOUND_WIDTH 1
`define I2C_I2C_STATUS_SLAVE_FOUND_LSB 0
`define I2C_I2C_STATUS_SLAVE_FOUND_MASK 32'h4
`define I2C_I2C_STATUS_SLAVE_FOUND_RESET 1'h0

// I2C_STATUS.TXE - Transmit register empty
`define I2C_I2C_STATUS_TXE_WIDTH 1
`define I2C_I2C_STATUS_TXE_LSB 1
`define I2C_I2C_STATUS_TXE_MASK 32'h4
`define I2C_I2C_STATUS_TXE_RESET 1'h1

// I2C_STATUS.TXNE - Transmit register not empty
`define I2C_I2C_STATUS_TXNE_WIDTH 1
`define I2C_I2C_STATUS_TXNE_LSB 2
`define I2C_I2C_STATUS_TXNE_MASK 32'h4
`define I2C_I2C_STATUS_TXNE_RESET 1'h0

// I2C_STATUS.RXE - Receive register empty
`define I2C_I2C_STATUS_RXE_WIDTH 1
`define I2C_I2C_STATUS_RXE_LSB 6
`define I2C_I2C_STATUS_RXE_MASK 32'h4
`define I2C_I2C_STATUS_RXE_RESET 1'h1

// I2C_STATUS.RXNE - Receive register not empty
`define I2C_I2C_STATUS_RXNE_WIDTH 1
`define I2C_I2C_STATUS_RXNE_LSB 7
`define I2C_I2C_STATUS_RXNE_MASK 32'h4
`define I2C_I2C_STATUS_RXNE_RESET 1'h0

// I2C_STATUS.ERR - Error flag
`define I2C_I2C_STATUS_ERR_WIDTH 1
`define I2C_I2C_STATUS_ERR_LSB 11
`define I2C_I2C_STATUS_ERR_MASK 32'h4
`define I2C_I2C_STATUS_ERR_RESET 1'h0

// I2C_STATUS.BUSY - I2C busy status
`define I2C_I2C_STATUS_BUSY_WIDTH 1
`define I2C_I2C_STATUS_BUSY_LSB 12
`define I2C_I2C_STATUS_BUSY_MASK 32'h4
`define I2C_I2C_STATUS_BUSY_RESET 1'h0

// I2C_STATUS.TS - Transmission complete
`define I2C_I2C_STATUS_TS_WIDTH 1
`define I2C_I2C_STATUS_TS_LSB 13
`define I2C_I2C_STATUS_TS_MASK 32'h4
`define I2C_I2C_STATUS_TS_RESET 1'h0

// I2C_STATUS.RS - Reception complete
`define I2C_I2C_STATUS_RS_WIDTH 1
`define I2C_I2C_STATUS_RS_LSB 14
`define I2C_I2C_STATUS_RS_MASK 32'h4
`define I2C_I2C_STATUS_RS_RESET 1'h0


// I2C_SLAVE_ADDR - I2C Slave Register Address
`define I2C_I2C_SLAVE_ADDR_ADDR 32'h8
`define I2C_I2C_SLAVE_ADDR_RESET 32'h0

// I2C_SLAVE_ADDR.ADDRESS - 8-bit register address
`define I2C_I2C_SLAVE_ADDR_ADDRESS_WIDTH 10
`define I2C_I2C_SLAVE_ADDR_ADDRESS_LSB 0
`define I2C_I2C_SLAVE_ADDR_ADDRESS_MASK 32'h8
`define I2C_I2C_SLAVE_ADDR_ADDRESS_RESET 10'h0


// I2C_REG_ADDR - I2C Slave Device Address
`define I2C_I2C_REG_ADDR_ADDR 32'hc
`define I2C_I2C_REG_ADDR_RESET 32'h0

// I2C_REG_ADDR.ADDS - 7 to 10-bit slave address
`define I2C_I2C_REG_ADDR_ADDS_WIDTH 8
`define I2C_I2C_REG_ADDR_ADDS_LSB 0
`define I2C_I2C_REG_ADDR_ADDS_MASK 32'hc
`define I2C_I2C_REG_ADDR_ADDS_RESET 8'h0


// I2C_TX_DATA_LOW - I2C Transmit Data Low 32-bit
`define I2C_I2C_TX_DATA_LOW_ADDR 32'h10
`define I2C_I2C_TX_DATA_LOW_RESET 32'h0

// I2C_TX_DATA_LOW.TX_DATA_LOW - Lower 32-bit of data to transmit
`define I2C_I2C_TX_DATA_LOW_TX_DATA_LOW_WIDTH 32
`define I2C_I2C_TX_DATA_LOW_TX_DATA_LOW_LSB 0
`define I2C_I2C_TX_DATA_LOW_TX_DATA_LOW_MASK 32'h10
`define I2C_I2C_TX_DATA_LOW_TX_DATA_LOW_RESET 32'h0


// I2C_TX_DATA_HIGH - I2C Transmit Data High 32-bit
`define I2C_I2C_TX_DATA_HIGH_ADDR 32'h14
`define I2C_I2C_TX_DATA_HIGH_RESET 32'h0

// I2C_TX_DATA_HIGH.TX_DATA_HIGH - Upper 32-bit of data to transmit
`define I2C_I2C_TX_DATA_HIGH_TX_DATA_HIGH_WIDTH 32
`define I2C_I2C_TX_DATA_HIGH_TX_DATA_HIGH_LSB 0
`define I2C_I2C_TX_DATA_HIGH_TX_DATA_HIGH_MASK 32'h14
`define I2C_I2C_TX_DATA_HIGH_TX_DATA_HIGH_RESET 32'h0


// I2C_RX_DATA_LOW - I2C Received Data Low 32-bit
`define I2C_I2C_RX_DATA_LOW_ADDR 32'h18
`define I2C_I2C_RX_DATA_LOW_RESET 32'h0

// I2C_RX_DATA_LOW.RX_DATA_LOW - Lower 32-bit of received data
`define I2C_I2C_RX_DATA_LOW_RX_DATA_LOW_WIDTH 32
`define I2C_I2C_RX_DATA_LOW_RX_DATA_LOW_LSB 0
`define I2C_I2C_RX_DATA_LOW_RX_DATA_LOW_MASK 32'h18
`define I2C_I2C_RX_DATA_LOW_RX_DATA_LOW_RESET 32'h0


// I2C_RX_DATA_HIGH - I2C Received Data High 32-bit
`define I2C_I2C_RX_DATA_HIGH_ADDR 32'h1c
`define I2C_I2C_RX_DATA_HIGH_RESET 32'h0

// I2C_RX_DATA_HIGH.RX_DATA_HIGH - Upper 32-bit of received data
`define I2C_I2C_RX_DATA_HIGH_RX_DATA_HIGH_WIDTH 32
`define I2C_I2C_RX_DATA_HIGH_RX_DATA_HIGH_LSB 0
`define I2C_I2C_RX_DATA_HIGH_RX_DATA_HIGH_MASK 32'h1c
`define I2C_I2C_RX_DATA_HIGH_RX_DATA_HIGH_RESET 32'h0


`endif // __REGS_I2C_VH