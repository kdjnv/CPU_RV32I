// Created with Corsair v1.0.4

`ifndef __REGS_GPIO_VH
`define __REGS_GPIO_VH

`define GPIO_BASE_ADDR 0
`define GPIO_DATA_WIDTH 32
`define GPIO_ADDR_WIDTH 32

// GPIO_IO - GPIO Read/Write Register
`define GPIO_GPIO_IO_ADDR 32'h0
`define GPIO_GPIO_IO_RESET 32'h0

// GPIO_IO.GPIO_0 - GPIO0
`define GPIO_GPIO_IO_GPIO_0_WIDTH 1
`define GPIO_GPIO_IO_GPIO_0_LSB 0
`define GPIO_GPIO_IO_GPIO_0_MASK 32'h0
`define GPIO_GPIO_IO_GPIO_0_RESET 1'h0

// GPIO_IO.GPIO_1 - GPIO1
`define GPIO_GPIO_IO_GPIO_1_WIDTH 1
`define GPIO_GPIO_IO_GPIO_1_LSB 1
`define GPIO_GPIO_IO_GPIO_1_MASK 32'h0
`define GPIO_GPIO_IO_GPIO_1_RESET 1'h0

// GPIO_IO.GPIO_2 - GPIO2
`define GPIO_GPIO_IO_GPIO_2_WIDTH 1
`define GPIO_GPIO_IO_GPIO_2_LSB 2
`define GPIO_GPIO_IO_GPIO_2_MASK 32'h0
`define GPIO_GPIO_IO_GPIO_2_RESET 1'h0

// GPIO_IO.GPIO_3 - GPIO3
`define GPIO_GPIO_IO_GPIO_3_WIDTH 1
`define GPIO_GPIO_IO_GPIO_3_LSB 3
`define GPIO_GPIO_IO_GPIO_3_MASK 32'h0
`define GPIO_GPIO_IO_GPIO_3_RESET 1'h0

// GPIO_IO.GPIO_4 - GPIO4
`define GPIO_GPIO_IO_GPIO_4_WIDTH 1
`define GPIO_GPIO_IO_GPIO_4_LSB 4
`define GPIO_GPIO_IO_GPIO_4_MASK 32'h0
`define GPIO_GPIO_IO_GPIO_4_RESET 1'h0

// GPIO_IO.GPIO_5 - GPIO5
`define GPIO_GPIO_IO_GPIO_5_WIDTH 1
`define GPIO_GPIO_IO_GPIO_5_LSB 5
`define GPIO_GPIO_IO_GPIO_5_MASK 32'h0
`define GPIO_GPIO_IO_GPIO_5_RESET 1'h0

// GPIO_IO.GPIO_6 - GPIO6
`define GPIO_GPIO_IO_GPIO_6_WIDTH 1
`define GPIO_GPIO_IO_GPIO_6_LSB 6
`define GPIO_GPIO_IO_GPIO_6_MASK 32'h0
`define GPIO_GPIO_IO_GPIO_6_RESET 1'h0

// GPIO_IO.GPIO_7 - GPIO7
`define GPIO_GPIO_IO_GPIO_7_WIDTH 1
`define GPIO_GPIO_IO_GPIO_7_LSB 7
`define GPIO_GPIO_IO_GPIO_7_MASK 32'h0
`define GPIO_GPIO_IO_GPIO_7_RESET 1'h0

// GPIO_IO.GPIO_8 - GPIO8
`define GPIO_GPIO_IO_GPIO_8_WIDTH 1
`define GPIO_GPIO_IO_GPIO_8_LSB 8
`define GPIO_GPIO_IO_GPIO_8_MASK 32'h0
`define GPIO_GPIO_IO_GPIO_8_RESET 1'h0

// GPIO_IO.GPIO_9 - GPIO9
`define GPIO_GPIO_IO_GPIO_9_WIDTH 1
`define GPIO_GPIO_IO_GPIO_9_LSB 9
`define GPIO_GPIO_IO_GPIO_9_MASK 32'h0
`define GPIO_GPIO_IO_GPIO_9_RESET 1'h0

// GPIO_IO.GPIO_10 - GPIO10
`define GPIO_GPIO_IO_GPIO_10_WIDTH 1
`define GPIO_GPIO_IO_GPIO_10_LSB 10
`define GPIO_GPIO_IO_GPIO_10_MASK 32'h0
`define GPIO_GPIO_IO_GPIO_10_RESET 1'h0

// GPIO_IO.GPIO_11 - GPIO11
`define GPIO_GPIO_IO_GPIO_11_WIDTH 1
`define GPIO_GPIO_IO_GPIO_11_LSB 11
`define GPIO_GPIO_IO_GPIO_11_MASK 32'h0
`define GPIO_GPIO_IO_GPIO_11_RESET 1'h0

// GPIO_IO.GPIO_12 - GPIO12
`define GPIO_GPIO_IO_GPIO_12_WIDTH 1
`define GPIO_GPIO_IO_GPIO_12_LSB 12
`define GPIO_GPIO_IO_GPIO_12_MASK 32'h0
`define GPIO_GPIO_IO_GPIO_12_RESET 1'h0

// GPIO_IO.GPIO_13 - GPIO13
`define GPIO_GPIO_IO_GPIO_13_WIDTH 1
`define GPIO_GPIO_IO_GPIO_13_LSB 13
`define GPIO_GPIO_IO_GPIO_13_MASK 32'h0
`define GPIO_GPIO_IO_GPIO_13_RESET 1'h0

// GPIO_IO.GPIO_14 - GPIO14
`define GPIO_GPIO_IO_GPIO_14_WIDTH 1
`define GPIO_GPIO_IO_GPIO_14_LSB 14
`define GPIO_GPIO_IO_GPIO_14_MASK 32'h0
`define GPIO_GPIO_IO_GPIO_14_RESET 1'h0

// GPIO_IO.GPIO_15 - GPIO15
`define GPIO_GPIO_IO_GPIO_15_WIDTH 1
`define GPIO_GPIO_IO_GPIO_15_LSB 15
`define GPIO_GPIO_IO_GPIO_15_MASK 32'h0
`define GPIO_GPIO_IO_GPIO_15_RESET 1'h0


// GPIO_CONFIG - GPIO_CONFIG
`define GPIO_GPIO_CONFIG_ADDR 32'h4
`define GPIO_GPIO_CONFIG_RESET 32'hff00

// GPIO_CONFIG.GPIO_0_CONFIG - GPIO0_CONFIG
`define GPIO_GPIO_CONFIG_GPIO_0_CONFIG_WIDTH 1
`define GPIO_GPIO_CONFIG_GPIO_0_CONFIG_LSB 0
`define GPIO_GPIO_CONFIG_GPIO_0_CONFIG_MASK 32'h4
`define GPIO_GPIO_CONFIG_GPIO_0_CONFIG_RESET 1'h0

// GPIO_CONFIG.GPIO_1_CONFIG - GPIO1_CONFIG
`define GPIO_GPIO_CONFIG_GPIO_1_CONFIG_WIDTH 1
`define GPIO_GPIO_CONFIG_GPIO_1_CONFIG_LSB 1
`define GPIO_GPIO_CONFIG_GPIO_1_CONFIG_MASK 32'h4
`define GPIO_GPIO_CONFIG_GPIO_1_CONFIG_RESET 1'h0

// GPIO_CONFIG.GPIO_2_CONFIG - GPIO2_CONFIG
`define GPIO_GPIO_CONFIG_GPIO_2_CONFIG_WIDTH 1
`define GPIO_GPIO_CONFIG_GPIO_2_CONFIG_LSB 2
`define GPIO_GPIO_CONFIG_GPIO_2_CONFIG_MASK 32'h4
`define GPIO_GPIO_CONFIG_GPIO_2_CONFIG_RESET 1'h0

// GPIO_CONFIG.GPIO_3_CONFIG - GPIO3_CONFIG
`define GPIO_GPIO_CONFIG_GPIO_3_CONFIG_WIDTH 1
`define GPIO_GPIO_CONFIG_GPIO_3_CONFIG_LSB 3
`define GPIO_GPIO_CONFIG_GPIO_3_CONFIG_MASK 32'h4
`define GPIO_GPIO_CONFIG_GPIO_3_CONFIG_RESET 1'h0

// GPIO_CONFIG.GPIO_4_CONFIG - GPIO4_CONFIG
`define GPIO_GPIO_CONFIG_GPIO_4_CONFIG_WIDTH 1
`define GPIO_GPIO_CONFIG_GPIO_4_CONFIG_LSB 4
`define GPIO_GPIO_CONFIG_GPIO_4_CONFIG_MASK 32'h4
`define GPIO_GPIO_CONFIG_GPIO_4_CONFIG_RESET 1'h0

// GPIO_CONFIG.GPIO_5_CONFIG - GPIO5_CONFIG
`define GPIO_GPIO_CONFIG_GPIO_5_CONFIG_WIDTH 1
`define GPIO_GPIO_CONFIG_GPIO_5_CONFIG_LSB 5
`define GPIO_GPIO_CONFIG_GPIO_5_CONFIG_MASK 32'h4
`define GPIO_GPIO_CONFIG_GPIO_5_CONFIG_RESET 1'h0

// GPIO_CONFIG.GPIO_6_CONFIG - GPIO6_CONFIG
`define GPIO_GPIO_CONFIG_GPIO_6_CONFIG_WIDTH 1
`define GPIO_GPIO_CONFIG_GPIO_6_CONFIG_LSB 6
`define GPIO_GPIO_CONFIG_GPIO_6_CONFIG_MASK 32'h4
`define GPIO_GPIO_CONFIG_GPIO_6_CONFIG_RESET 1'h0

// GPIO_CONFIG.GPIO_7_CONFIG - GPIO7_CONFIG
`define GPIO_GPIO_CONFIG_GPIO_7_CONFIG_WIDTH 1
`define GPIO_GPIO_CONFIG_GPIO_7_CONFIG_LSB 7
`define GPIO_GPIO_CONFIG_GPIO_7_CONFIG_MASK 32'h4
`define GPIO_GPIO_CONFIG_GPIO_7_CONFIG_RESET 1'h0

// GPIO_CONFIG.GPIO_8_CONFIG - GPIO8_CONFIG
`define GPIO_GPIO_CONFIG_GPIO_8_CONFIG_WIDTH 1
`define GPIO_GPIO_CONFIG_GPIO_8_CONFIG_LSB 8
`define GPIO_GPIO_CONFIG_GPIO_8_CONFIG_MASK 32'h4
`define GPIO_GPIO_CONFIG_GPIO_8_CONFIG_RESET 1'h1

// GPIO_CONFIG.GPIO_9_CONFIG - GPIO9_CONFIG
`define GPIO_GPIO_CONFIG_GPIO_9_CONFIG_WIDTH 1
`define GPIO_GPIO_CONFIG_GPIO_9_CONFIG_LSB 9
`define GPIO_GPIO_CONFIG_GPIO_9_CONFIG_MASK 32'h4
`define GPIO_GPIO_CONFIG_GPIO_9_CONFIG_RESET 1'h1

// GPIO_CONFIG.GPIO_10_CONFIG - GPIO10_CONFIG
`define GPIO_GPIO_CONFIG_GPIO_10_CONFIG_WIDTH 1
`define GPIO_GPIO_CONFIG_GPIO_10_CONFIG_LSB 10
`define GPIO_GPIO_CONFIG_GPIO_10_CONFIG_MASK 32'h4
`define GPIO_GPIO_CONFIG_GPIO_10_CONFIG_RESET 1'h1

// GPIO_CONFIG.GPIO_11_CONFIG - GPIO11_CONFIG
`define GPIO_GPIO_CONFIG_GPIO_11_CONFIG_WIDTH 1
`define GPIO_GPIO_CONFIG_GPIO_11_CONFIG_LSB 11
`define GPIO_GPIO_CONFIG_GPIO_11_CONFIG_MASK 32'h4
`define GPIO_GPIO_CONFIG_GPIO_11_CONFIG_RESET 1'h1

// GPIO_CONFIG.GPIO_12_CONFIG - GPIO12_CONFIG
`define GPIO_GPIO_CONFIG_GPIO_12_CONFIG_WIDTH 1
`define GPIO_GPIO_CONFIG_GPIO_12_CONFIG_LSB 12
`define GPIO_GPIO_CONFIG_GPIO_12_CONFIG_MASK 32'h4
`define GPIO_GPIO_CONFIG_GPIO_12_CONFIG_RESET 1'h1

// GPIO_CONFIG.GPIO_13_CONFIG - GPIO13_CONFIG
`define GPIO_GPIO_CONFIG_GPIO_13_CONFIG_WIDTH 1
`define GPIO_GPIO_CONFIG_GPIO_13_CONFIG_LSB 13
`define GPIO_GPIO_CONFIG_GPIO_13_CONFIG_MASK 32'h4
`define GPIO_GPIO_CONFIG_GPIO_13_CONFIG_RESET 1'h1

// GPIO_CONFIG.GPIO_14_CONFIG - GPIO14_CONFIG
`define GPIO_GPIO_CONFIG_GPIO_14_CONFIG_WIDTH 1
`define GPIO_GPIO_CONFIG_GPIO_14_CONFIG_LSB 14
`define GPIO_GPIO_CONFIG_GPIO_14_CONFIG_MASK 32'h4
`define GPIO_GPIO_CONFIG_GPIO_14_CONFIG_RESET 1'h1

// GPIO_CONFIG.GPIO_15_CONFIG - GPIO15_CONFIG
`define GPIO_GPIO_CONFIG_GPIO_15_CONFIG_WIDTH 1
`define GPIO_GPIO_CONFIG_GPIO_15_CONFIG_LSB 15
`define GPIO_GPIO_CONFIG_GPIO_15_CONFIG_MASK 32'h4
`define GPIO_GPIO_CONFIG_GPIO_15_CONFIG_RESET 1'h1


`endif // __REGS_GPIO_VH